// Copyright 2016-2024 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


parameter vpiFunction = 20;
parameter vpiIODecl = 28;
parameter vpiModule = 32;
parameter vpiParameter = 41;
parameter vpiTask = 59;

parameter vpiAttribute = 105;

parameter vpiExpr = 102;
parameter vpiFrame = 110;

parameter vpiPackage = 600;
parameter vpiTypespec = 605;

parameter vpiStringVar = 616;

parameter vpiIntTypespec = 629;
parameter vpiClassTypespec = 630;

parameter vpiClassDefn = 652;
parameter vpiExtends = 677;
