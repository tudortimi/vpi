module some_module #(
    parameter bit SOME_BIT_PARAM = 0,
    parameter int SOME_INT_PARAM = 42);
endmodule
