// Copyright 2016-2024 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


parameter vpiLhs = 77;
parameter vpiRhs = 82;
parameter vpiScope = 84;

parameter vpiClassObj = 621;

parameter vpiReturn = 666;
parameter vpiOrigin = 713;
parameter vpiPrefix = 714;
parameter vpiInstance = 745;
