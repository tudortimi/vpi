// Copyright 2016 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


parameter vpiUndefined = -1;
parameter vpiType = 1;
parameter vpiName = 2;
parameter vpiFullName = 3;
parameter vpiDefName = 9;
parameter vpiTimeUnit = 11;
parameter vpiTimePrecision = 12;

parameter vpiDirection = 20;
parameter vpiInput = 1;
parameter vpiOutput = 2;
parameter vpiInout = 3;

parameter vpiActive = 49;
parameter vpiAutomatic = 50;
parameter vpiConstantVariable = 612;

parameter vpiRandType = 610;
parameter vpiNotRand = 1;
parameter vpiRand = 2;
parameter vpiRandC = 3;

parameter vpiVirtual = 635;

parameter vpiMethod = 645;
parameter vpiObjId = 660;
