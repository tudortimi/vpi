module some_module #(
    parameter bit SOME_BIT_PARAM = 0,
    parameter int SOME_INT_PARAM = 42,
    parameter int SOME_OTHER_INT_PARAM = 1000);
endmodule
